`define DELAY 30
module _alu_testbench();

reg [31:0] a;
reg [31:0] b;
reg [2:0] opCode;
wire [31:0] result;
wire ZERO;

alu32 al(result,ZERO,a,b,opCode);

initial begin

opCode = 3'b000;
a = 32'b00000010101010001100111111111111;
b = 32'b11111000000000000000000000111111;
#`DELAY
opCode = 3'b000;
a = 32'b00000010101010001100111111111111;
b = 32'b00000010101010001100111111111111;
#`DELAY
opCode = 3'b000;
a = 32'b00000000000000000000111111111111;
b = 32'b11111111111111111111110000000000;
/////////////////////////////////////////
#`DELAY
opCode = 3'b001;
a = 32'b11111111111111111111111111111111;
b = 32'b00000000000000000000000000000000;
#`DELAY
opCode = 3'b001;
a = 32'b10101010101010101010101010101010;
b = 32'b01010101010101010101010101010101;
#`DELAY
opCode = 3'b001;
a = 32'b01010000000000001011111111111111;
b = 32'b00000000000000000000011111111111;
/////////////////////////////////////////
#`DELAY
opCode = 3'b010;
a = 32'b00000000000000000000000000000000;
b = 32'b11111111111111111111111111111111;
#`DELAY
opCode = 3'b010;
a = 32'b00111111111111111111111111111111;
b = 32'b00111111111111111111111111111111;
#`DELAY
opCode = 3'b010;
a = 32'b00000000000000000000000000011111;
b = 32'b00000000000000000000000000011111;
/////////////////////////////////////////
#`DELAY
opCode = 3'b011;
a = 32'b11111111111111111111111111111111;
b = 32'b00000000000000000000000000000000;
#`DELAY
opCode = 3'b011;
a = 32'b11111111111111111111111111111111;
b = 32'b11111111111111111111111111111111;
#`DELAY
opCode = 3'b011;
a = 32'b10101010101010101010101010101010;
b = 32'b01010101010101010101010101010101;
/////////////////////////////////////////
#`DELAY
opCode = 3'b100;
a = 32'b10000111111111111111111111111111;
b = 32'b10000111111111111111111111111111;
#`DELAY
opCode = 3'b100;
a = 32'b00000000000000000111111111111111;
b = 32'b00000000000000000000000000001111;
#`DELAY
opCode = 3'b100;
a = 32'b00000000000000000000000000011111;
b = 32'b00000000000000000000000000000000;
/////////////////////////////////////////
#`DELAY
opCode = 3'b101;
a = 32'b10000000000000000111111111111111;
b = 32'b00000000000000000000000000000011;
#`DELAY
opCode = 3'b101;
a = 32'b10000000000000000000000000000000;
b = 32'b00000000000000000000000000011111;
#`DELAY
opCode = 3'b101;
a = 32'b11111111111111111111111111111111;
b = 32'b00000000000000000000000100000000;
/////////////////////////////////////////
#`DELAY
opCode = 3'b110;
a = 32'b11111111111111111111111111111111;
b = 32'b00000000000000000000000000000100;
#`DELAY
opCode = 3'b110;
a = 32'b00000000000000011111111111111111;
b = 32'b00000000000000000000000000001111;
#`DELAY
opCode = 3'b110;
a = 32'b11111111111111111111111111111111;
b = 32'b00000000000000011111000010000000;
/////////////////////////////////////////
#`DELAY
opCode = 3'b111;
a = 32'b11111111111111111111111111111111;
b = 32'b00000000000000000000000000000000;
#`DELAY
opCode = 3'b111;
a = 32'b00000000000000111111111111111111;
b = 32'b00000000000000111111111111111111;
#`DELAY
opCode = 3'b111;
a = 32'b10101010101010101010101010101010;
b = 32'b00000000000000000000000000000000;
/////////////////////////////////////////



end

initial begin

$monitor("a = %32b , b = %32b ,OPCODE = %3b ,result = %32b ,ZERO = %1b",a,b,opCode,result,ZERO);
end
endmodule